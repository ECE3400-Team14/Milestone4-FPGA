`define SCREEN_WIDTH 176
`define SCREEN_HEIGHT 144

///////* DON'T CHANGE THIS PART *///////
module DE0_NANO(
	CLOCK_50,
	GPIO_0_D,
	GPIO_1_D,
	KEY,
	LED
);

//=======================================================
//  PARAMETER declarations
//=======================================================
localparam RED = 8'b111_000_00;
localparam GREEN = 8'b000_111_00;
localparam BLUE = 8'b000_000_11;

//=======================================================
//  PORT declarations
//=======================================================

//////////// CLOCK - DON'T NEED TO CHANGE THIS //////////
input 		          		CLOCK_50;

//////////// GPIO_0, GPIO_0 connect to GPIO Default //////////
output 		    [33:0]		GPIO_0_D;
output          [7:0]      LED;
//////////// GPIO_0, GPIO_1 connect to GPIO Default //////////
input 		    [33:0]		GPIO_1_D;
input 		     [1:0]		KEY;

///// PIXEL DATA /////
wire [7:0]	pixel_data_RGB332;

///// READ/WRITE ADDRESS /////
wire [14:0] X_ADDR;
wire [14:0] Y_ADDR;
wire [14:0] WRITE_ADDRESS;
reg [14:0] READ_ADDRESS; 

assign WRITE_ADDRESS = X_ADDR + Y_ADDR*(`SCREEN_WIDTH);

///// VGA INPUTS/OUTPUTS /////
wire 			VGA_RESET;
wire [7:0]	VGA_COLOR_IN;
wire [9:0]	VGA_PIXEL_X;
wire [9:0]	VGA_PIXEL_Y;
wire [7:0]	MEM_OUTPUT;
wire			VGA_VSYNC_NEG;
wire			VGA_HSYNC_NEG;
reg			VGA_READ_MEM_EN;

assign GPIO_0_D[5] = VGA_VSYNC_NEG;
assign GPIO_0_D[31] = c0_sig;
assign VGA_RESET = ~KEY[0];

///// I/O for Img Proc /////
wire [8:0] RESULT;

/* WRITE ENABLE */
wire W_EN;

///////* CREATE ANY LOCAL WIRES YOU NEED FOR YOUR PLL *///////
wire c0_sig;
wire c1_sig;
wire c2_sig;

//SIM
wire VSYNC;
wire HREF;
wire [7:0] sim_data;

///////* INSTANTIATE YOUR PLL HERE *///////

PLL	PLL_inst (
	.inclk0 ( CLOCK_50 ),
	.c0 ( c0_sig ),
	.c1 ( c1_sig ),
	.c2 ( c2_sig )
	);

///////* M9K Module *///////
Dual_Port_RAM_M9K mem(
	.input_data(pixel_data_RGB332),
	.w_addr(WRITE_ADDRESS),
	.r_addr(READ_ADDRESS),
	.w_en(W_EN),
	.clk_W(c2_sig),
	.clk_R(c1_sig), // DO WE NEED TO READ SLOWER THAN WRITE??
	.output_data(MEM_OUTPUT)
);

///////* VGA Module *///////
VGA_DRIVER driver (
	.RESET(VGA_RESET),
	.CLOCK(c1_sig),
	.PIXEL_COLOR_IN(VGA_READ_MEM_EN ? MEM_OUTPUT : BLUE),
	.PIXEL_X(VGA_PIXEL_X),
	.PIXEL_Y(VGA_PIXEL_Y),
	.PIXEL_COLOR_OUT({GPIO_0_D[9],GPIO_0_D[11],GPIO_0_D[13],GPIO_0_D[15],GPIO_0_D[17],GPIO_0_D[19],GPIO_0_D[21],GPIO_0_D[23]}),
   .H_SYNC_NEG(GPIO_0_D[7]),
   .V_SYNC_NEG(VGA_VSYNC_NEG)
);

///////* Image Processor *///////
IMAGE_PROCESSOR proc(
	.PIXEL_IN(MEM_OUTPUT),
	.CLK(c1_sig),
	.VGA_PIXEL_X(VGA_PIXEL_X),
	.VGA_PIXEL_Y(VGA_PIXEL_Y),
	.VGA_VSYNC_NEG(VGA_VSYNC_NEG),
	.RESULT(RESULT),
	.shape(shape),
	.top(),
	.bottom(),
	.first(),
	.second(),
	.third(),
	.colorFinished(colorFinished),
	.shapeFinished(shapeFinished),
	.red(),
	.blue(red)
);
wire [14:0] red;
wire [1:0] shape;
//assign LED = red[7:0];
//assign LED = {2'b0,shape, RESULT[1],RESULT[1],RESULT[0],RESULT[0]};

//communicate to Arduino
SERIAL serial(
	.CLK(c1_sig),
	.RESULT(RESULT),
	.colorFinished(colorFinished),
	.shapeFinished(shapeFinished),
	.shape(shape),
	.SIG(GPIO_1_D[32]),
	.DATA(GPIO_0_D[33]),
	.write(write),
	.SHAPE_DATA(LED)
);
wire colorFinished;
wire shapeFinished;
wire [3:0] write;
//assign LED = {write};//, GPIO_1_D[32],GPIO_0_D[33]};

//
//SIMULATOR simulator(
//  .CLK(c0_sig),
//  .VSYNC(VSYNC),
//  .HREF(HREF),
//  .DATA(sim_data)
//);

SIMULATOR_OLD simulator(
  .CLK(c0_sig),
  .VSYNC(VSYNC),
  .HREF(HREF),
  .DATA(sim_data)
);

 
// simulator control unit
//CONTROL_UNIT control_unit(
//  .CLK(c0_sig),
//  .HREF(HREF),
//  .VSYNC(VSYNC),
//  .input_data(sim_data),
//  .output_data(pixel_data_RGB332),
//  .X_ADDR(X_ADDR),
//  .Y_ADDR(Y_ADDR),
//  .w_en(W_EN)
//);

//camera control unit
CONTROL_UNIT control_unit(
  .CLK(GPIO_1_D[13]),
  .HREF(GPIO_1_D[15]),
  .VSYNC(GPIO_1_D[14]),
  .input_data(GPIO_1_D[23:16]),
  .output_data(pixel_data_RGB332),
  .X_ADDR(X_ADDR),
  .Y_ADDR(Y_ADDR),
  .w_en(W_EN)
);

///////* Update Read Address *///////
always @ (VGA_PIXEL_X, VGA_PIXEL_Y) begin
		READ_ADDRESS = (VGA_PIXEL_X + VGA_PIXEL_Y*`SCREEN_WIDTH);
		if(VGA_PIXEL_X>(`SCREEN_WIDTH-1) || VGA_PIXEL_Y>(`SCREEN_HEIGHT-1)) begin
				VGA_READ_MEM_EN = 1'b0;
		end
		else begin
				VGA_READ_MEM_EN = 1'b1;
		end
end
//wire [7:0] part;
//assign LED[7:0] = GPIO_1_D[23:16];
//assign LED[7:4] = shape;
//assign LED[3:0] = RESULT[3:0];
//assign LED[0] = pixel_data_RGB332[7];
//assign LED[1] = pixel_data_RGB332[6];
//assign LED[2] = pixel_data_RGB332[5];
//assign LED[3] = pixel_data_RGB332[4];
//assign LED[4] = pixel_data_RGB332[3];
//assign LED[5] = pixel_data_RGB332[2];
//assign LED[6] = pixel_data_RGB332[1];
//assign LED[7] = pixel_data_RGB332[0];
	
endmodule 